--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   06:48:33 04/15/2024
-- Design Name:   
-- Module Name:   D:/Student/Desktop/NADAABOSAADA 211002838/datamemtest.vhd
-- Project Name:  mips211002838nadafouadfinal
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: DataMemory
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY datamemtest IS
END datamemtest;
 
ARCHITECTURE behavior OF datamemtest IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT DataMemory
    PORT(
         Address : IN  std_logic_vector(31 downto 0);
         readdata : OUT  std_logic_vector(31 downto 0);
         writedata : IN  std_logic_vector(31 downto 0);
         clk : IN  std_logic;
         memread : IN  std_logic;
         memwrite : IN  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal Address : std_logic_vector(31 downto 0) := (others => '0');
   signal writedata : std_logic_vector(31 downto 0) := (others => '0');
   signal clk : std_logic := '0';
   signal memread : std_logic := '0';
   signal memwrite : std_logic := '0';

 	--Outputs
   signal readdata : std_logic_vector(31 downto 0);

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: DataMemory PORT MAP (
          Address => Address,
          readdata => readdata,
          writedata => writedata,
          clk => clk,
          memread => memread,
          memwrite => memwrite
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
		
		
      wait for 100 ns;	

      wait for clk_period*10;

      -- insert stimulus here
		memread>='0';	
		memwrite>='1';
		Address>= X"00000000";
		writedata>= "00001111000011110000111100001111";
		
		wait for 100 ns;
		
		memread>='1';	
		memwrite>='0';
		Address>= X"00000001";
		wait for 100 ns;

      wait;
   end process;

END;
